module risc_v_core (
  input
  output
);

endmodule
