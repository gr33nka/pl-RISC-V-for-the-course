module hazard_unit (
  input 
  output
);


endmodule
