module writeback (
  input       [ : ] ,
  output  reg [ : ] ,
);

endmodule
