module memory (
  input       [ : ] ,
  output  reg [ : ] ,
);

endmodule
