module execute (
  input       [ : ] ,
  output  reg [ : ] ,
);

endmodule
