module decode (
  input       [ : ] ,
  output  reg [ : ] ,
);

endmodule
