module fetch (
  input       [ : ] ,
  output  reg [ : ] ,
);

endmodule
